library verilog;
use verilog.vl_types.all;
entity \topic__2_1_vlg_vec_tst\ is
end \topic__2_1_vlg_vec_tst\;
