library verilog;
use verilog.vl_types.all;
entity \topic__2_3\ is
    port(
        \Out\           : out    vl_logic;
        F               : in     vl_logic;
        E               : in     vl_logic;
        G               : in     vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic
    );
end \topic__2_3\;
