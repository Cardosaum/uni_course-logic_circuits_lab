library verilog;
use verilog.vl_types.all;
entity \topic__2_3_vlg_check_tst\ is
    port(
        \Out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end \topic__2_3_vlg_check_tst\;
